module cmp 
(
    clk,reset,inst_in,d_in,pc_out,d_out,addr_out,memWrEn,memEn
);
    
endmodule