module ID (
    clk,reset,ID_inst,ID_pc,
    ID_flush
);
    input wire clk,reset;
    input wire [0:31] ID_inst, ID_pc;

    output ID_flush;
    //branch and hdu

    


endmodule